module test
    or
    and
    xor
endmodule